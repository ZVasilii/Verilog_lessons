module top(input CLK);

endmodule